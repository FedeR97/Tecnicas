-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
-- CREATED		"Fri Oct 24 21:17:01 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

	PORT
	(
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		A2 :  IN  STD_LOGIC;
		A3 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		P0 :  OUT  STD_LOGIC;
		P1 :  OUT  STD_LOGIC;
		P2 :  OUT  STD_LOGIC;
		P3 :  OUT  STD_LOGIC;
		P4 :  OUT  STD_LOGIC;
		P5 :  OUT  STD_LOGIC;
		P6 :  OUT  STD_LOGIC;
		P7 :  OUT  STD_LOGIC
	);
END MultiB;

ARCHITECTURE bdf_type OF MultiB IS 

COMPONENT sumador_completo
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CI : IN STD_LOGIC;
		 CO : OUT STD_LOGIC;
		 S : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	A0C :  STD_LOGIC;
SIGNAL	A1C :  STD_LOGIC;
SIGNAL	A2C :  STD_LOGIC;
SIGNAL	A3C :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_2 <= '0';
SYNTHESIZED_WIRE_14 <= '0';
SYNTHESIZED_WIRE_22 <= '0';
SYNTHESIZED_WIRE_26 <= '0';



SYNTHESIZED_WIRE_13 <= B1 AND A0C;


b2v_inst10 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_1,
		 CI => SYNTHESIZED_WIRE_2,
		 CO => SYNTHESIZED_WIRE_5,
		 S => P3);


b2v_inst11 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_3,
		 B => SYNTHESIZED_WIRE_4,
		 CI => SYNTHESIZED_WIRE_5,
		 CO => SYNTHESIZED_WIRE_8,
		 S => P4);


b2v_inst12 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_6,
		 B => SYNTHESIZED_WIRE_7,
		 CI => SYNTHESIZED_WIRE_8,
		 CO => SYNTHESIZED_WIRE_11,
		 S => P5);


b2v_inst13 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_9,
		 B => SYNTHESIZED_WIRE_10,
		 CI => SYNTHESIZED_WIRE_11,
		 CO => P7,
		 S => P6);


P0 <= B0 AND A0C;


SYNTHESIZED_WIRE_12 <= B0 AND A1C;



SYNTHESIZED_WIRE_16 <= B0 AND A2C;


SYNTHESIZED_WIRE_19 <= B0 AND A3C;


SYNTHESIZED_WIRE_15 <= B1 AND A1C;


b2v_inst2 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_12,
		 B => SYNTHESIZED_WIRE_13,
		 CI => SYNTHESIZED_WIRE_14,
		 CO => SYNTHESIZED_WIRE_17,
		 S => P1);


SYNTHESIZED_WIRE_18 <= B1 AND A2C;


SYNTHESIZED_WIRE_21 <= B1 AND A3C;



SYNTHESIZED_WIRE_24 <= B2 AND A0C;


SYNTHESIZED_WIRE_27 <= B2 AND A1C;


SYNTHESIZED_WIRE_30 <= B2 AND A2C;


SYNTHESIZED_WIRE_33 <= B2 AND A3C;


SYNTHESIZED_WIRE_0 <= B3 AND A0C;


SYNTHESIZED_WIRE_3 <= B3 AND A1C;


SYNTHESIZED_WIRE_6 <= B3 AND A2C;


b2v_inst3 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_15,
		 B => SYNTHESIZED_WIRE_16,
		 CI => SYNTHESIZED_WIRE_17,
		 CO => SYNTHESIZED_WIRE_20,
		 S => SYNTHESIZED_WIRE_25);


SYNTHESIZED_WIRE_9 <= B3 AND A3C;




b2v_inst4 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_18,
		 B => SYNTHESIZED_WIRE_19,
		 CI => SYNTHESIZED_WIRE_20,
		 CO => SYNTHESIZED_WIRE_23,
		 S => SYNTHESIZED_WIRE_28);


b2v_inst5 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_21,
		 B => SYNTHESIZED_WIRE_22,
		 CI => SYNTHESIZED_WIRE_23,
		 CO => SYNTHESIZED_WIRE_34,
		 S => SYNTHESIZED_WIRE_31);


b2v_inst6 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_24,
		 B => SYNTHESIZED_WIRE_25,
		 CI => SYNTHESIZED_WIRE_26,
		 CO => SYNTHESIZED_WIRE_29,
		 S => P2);


b2v_inst7 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_27,
		 B => SYNTHESIZED_WIRE_28,
		 CI => SYNTHESIZED_WIRE_29,
		 CO => SYNTHESIZED_WIRE_32,
		 S => SYNTHESIZED_WIRE_1);


b2v_inst8 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_30,
		 B => SYNTHESIZED_WIRE_31,
		 CI => SYNTHESIZED_WIRE_32,
		 CO => SYNTHESIZED_WIRE_35,
		 S => SYNTHESIZED_WIRE_4);


b2v_inst9 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_33,
		 B => SYNTHESIZED_WIRE_34,
		 CI => SYNTHESIZED_WIRE_35,
		 CO => SYNTHESIZED_WIRE_10,
		 S => SYNTHESIZED_WIRE_7);

A0C <= A0;
A1C <= A1;
A2C <= A2;
A3C <= A3;

END bdf_type;