-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Thu Oct 30 23:26:04 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ParteE IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        z1 : OUT STD_LOGIC;
        z2 : OUT STD_LOGIC;
        z3 : OUT STD_LOGIC;
        z4 : OUT STD_LOGIC;
        z5 : OUT STD_LOGIC;
        z6 : OUT STD_LOGIC;
        z7 : OUT STD_LOGIC
    );
END ParteE;

ARCHITECTURE BEHAVIOR OF ParteE IS
    TYPE type_fstate IS (state4,state2,state3,state7,state6,state5,state1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            z1 <= '0';
            z2 <= '0';
            z3 <= '0';
            z4 <= '0';
            z5 <= '0';
            z6 <= '0';
            z7 <= '0';
        ELSE
            z1 <= '0';
            z2 <= '0';
            z3 <= '0';
            z4 <= '0';
            z5 <= '0';
            z6 <= '0';
            z7 <= '0';
            CASE fstate IS
                WHEN state4 =>
                    reg_fstate <= state1;

                    z4 <= '1';
                WHEN state2 =>
                    reg_fstate <= state3;

                    z2 <= '1';
                WHEN state3 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= state4;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    z3 <= '1';
                WHEN state7 =>
                    reg_fstate <= state1;

                    z7 <= '1';
                WHEN state6 =>
                    reg_fstate <= state3;

                    z6 <= '1';
                WHEN state5 =>
                    reg_fstate <= state6;

                    z5 <= '1';
                WHEN state1 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= state2;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    z1 <= '1';
                WHEN OTHERS => 
                    z1 <= 'X';
                    z2 <= 'X';
                    z3 <= 'X';
                    z4 <= 'X';
                    z5 <= 'X';
                    z6 <= 'X';
                    z7 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
