-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Fri Oct 31 11:13:01 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY I2Control IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SDA : IN STD_LOGIC := '0';
        SOY : IN STD_LOGIC := '0';
        Fin_dato : IN STD_LOGIC := '0';
        Fin_dir : IN STD_LOGIC := '0';
        Hab_dir : OUT STD_LOGIC;
        Hab_dato : OUT STD_LOGIC
    );
END I2Control;

ARCHITECTURE BEHAVIOR OF I2Control IS
    TYPE type_fstate IS (Oscioso,Guardar_Dir,R_W,ACK,Guardar_dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,SOY,Fin_dato,Fin_dir)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            Hab_dir <= '0';
            Hab_dato <= '0';
        ELSE
            Hab_dir <= '0';
            Hab_dato <= '0';
            CASE fstate IS
                WHEN Oscioso =>
                    IF ((SDA = '0')) THEN
                        reg_fstate <= Guardar_Dir;
                    ELSIF ((SDA = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    Hab_dato <= '0';

                    Hab_dir <= '0';
                WHEN Guardar_Dir =>
                    IF (((Fin_dir = '1') AND (SOY = '1'))) THEN
                        reg_fstate <= R_W;
                    ELSIF ((Fin_dir = '0')) THEN
                        reg_fstate <= Guardar_Dir;
                    ELSIF (((Fin_dir = '1') AND (SOY = '0'))) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_Dir;
                    END IF;

                    Hab_dato <= '0';

                    Hab_dir <= '1';
                WHEN R_W =>
                    reg_fstate <= ACK;

                    Hab_dato <= '0';

                    Hab_dir <= '0';
                WHEN ACK =>
                    reg_fstate <= Guardar_dato;

                    Hab_dato <= '0';

                    Hab_dir <= '0';
                WHEN Guardar_dato =>
                    IF ((Fin_dato = '0')) THEN
                        reg_fstate <= Guardar_dato;
                    ELSIF ((Fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_dato;
                    END IF;

                    Hab_dato <= '1';

                    Hab_dir <= '0';
                WHEN OTHERS => 
                    Hab_dir <= 'X';
                    Hab_dato <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
